/*
 * Microgreen Growth Classifier - TinyTapeout tt08
 * 
 * AI-powered growth stage detection for precision farming
 * Training accuracy: 89.4% | Test accuracy: 86.7%
 * 
 * Classes: 0 = Not Ready (Growing), 1 = Ready to Harvest
 * Architecture: 4 inputs → 4 hidden neurons → 2 outputs
 */

module tt_um_microgreen_classifier (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (bidirectional)
    input  wire       ena,      // Enable - will go high when design is enabled
    input  wire       clk,      // Clock - 50MHz
    input  wire       rst_n     // Reset - active low
);

    // Configure all bidirectional pins as outputs
    assign uio_oe = 8'b11111111;
    assign uio_out = 8'b00000000;  // Not used in this version

    // ========================================================================
    // INPUT PIN MAPPING
    // ========================================================================
    // ui_in[3:0] - Height sensor (4 bits, 0-15 scale)
    // ui_in[7:4] - Color/Greenness sensor (4 bits, 0-15 scale)
    // uio_in[3:0] - Density sensor (4 bits, 0-15 scale)
    // uio_in[7:4] - Texture/Temperature sensor (4 bits, 0-15 scale)
    
    wire [3:0] feature_height = ui_in[3:0];
    wire [3:0] feature_color = ui_in[7:4];
    wire [3:0] feature_density = uio_in[3:0];
    wire [3:0] feature_texture = uio_in[7:4];

    // ========================================================================
    // TRAINED WEIGHTS - UPDATE THESE FROM weights.vh
    // ========================================================================
    // TODO: Open your weights.vh file and copy the parameter values here!
    // These are PLACEHOLDER values - replace with YOUR trained weights
    
    // Input to Hidden Layer Weights (4 neurons × 4 inputs)
    parameter [3:0] W_IH_0 = 4'b1001;  // REPLACE with your W_IH_0
    parameter [3:0] W_IH_1 = 4'b1011;  // REPLACE with your W_IH_1
    parameter [3:0] W_IH_2 = 4'b1100;  // REPLACE with your W_IH_2
    parameter [3:0] W_IH_3 = 4'b1110;  // REPLACE with your W_IH_3
    
    // Hidden to Output Layer Weights (2 neurons × 4 hidden)
    parameter [3:0] W_HO_0 = 4'b1010;  // REPLACE with your W_HO_0
    parameter [3:0] W_HO_1 = 4'b0101;  // REPLACE with your W_HO_1
    
    // Hidden Layer Biases
    parameter signed [3:0] BIAS_H0 = 4'sd1;  // REPLACE with your BIAS_H0
    parameter signed [3:0] BIAS_H1 = 4'sd1;  // REPLACE with your BIAS_H1
    parameter signed [3:0] BIAS_H2 = -4'sd1;  // REPLACE with your BIAS_H2
    parameter signed [3:0] BIAS_H3 = 4'sd1;  // REPLACE with your BIAS_H3

    // ========================================================================
    // STATE MACHINE
    // ========================================================================
    reg [2:0] state;
    localparam IDLE = 3'd0;
    localparam COMPUTE_HIDDEN = 3'd1;
    localparam COMPUTE_OUTPUT = 3'd2;
    localparam DONE = 3'd3;
    
    // Registers
    reg [3:0] hidden_act;      // Hidden layer activations
    reg classification;         // Output: 0=not ready, 1=ready
    reg ready;                 // Result ready flag
    
    // ========================================================================
    // XNOR-POPCOUNT FUNCTION (Core BNN Operation)
    // ========================================================================
    function [4:0] xnor_popcount;
        input [3:0] a;
        input [3:0] b;
        reg [3:0] xnor_result;
        integer i, count;
        begin
            xnor_result = ~(a ^ b);  // XNOR: 1 when bits match
            count = 0;
            for (i = 0; i < 4; i = i + 1) begin
                if (xnor_result[i]) count = count + 1;
            end
            xnor_popcount = count;
        end
    endfunction
    
    // ========================================================================
    // BINARIZATION FUNCTION
    // ========================================================================
    function binarize;
        input [3:0] val;
        begin
            binarize = (val >= 4'd8) ? 1'b1 : 1'b0;  // Threshold at midpoint
        end
    endfunction
    
    // ========================================================================
    // LAYER 1: HIDDEN LAYER COMPUTATION
    // ========================================================================
    
    // Binarize all inputs
    wire [3:0] inputs_binary = {
        binarize(feature_texture),
        binarize(feature_density),
        binarize(feature_color),
        binarize(feature_height)
    };
    
    // Compute weighted sums for hidden neurons
    wire signed [4:0] hidden_sum [0:3];
    assign hidden_sum[0] = xnor_popcount(inputs_binary, W_IH_0) + BIAS_H0 - 2;
    assign hidden_sum[1] = xnor_popcount(inputs_binary, W_IH_1) + BIAS_H1 - 2;
    assign hidden_sum[2] = xnor_popcount(inputs_binary, W_IH_2) + BIAS_H2 - 2;
    assign hidden_sum[3] = xnor_popcount(inputs_binary, W_IH_3) + BIAS_H3 - 2;
    
    // ========================================================================
    // LAYER 2: OUTPUT LAYER COMPUTATION
    // ========================================================================
    
    // Compute output scores
    wire signed [4:0] output_sum [0:1];
    assign output_sum[0] = xnor_popcount(hidden_act, W_HO_0);  // Score for "not ready"
    assign output_sum[1] = xnor_popcount(hidden_act, W_HO_1);  // Score for "ready"
    
    // Winner-take-all decision
    wire decision = (output_sum[1] > output_sum[0]) ? 1'b1 : 1'b0;
    
    // ========================================================================
    // STATE MACHINE LOGIC
    // ========================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= IDLE;
            hidden_act <= 4'b0;
            classification <= 1'b0;
            ready <= 1'b0;
        end else if (ena) begin
            case (state)
                IDLE: begin
                    ready <= 1'b0;
                    state <= COMPUTE_HIDDEN;
                end
                
                COMPUTE_HIDDEN: begin
                    // Apply sign activation function
                    hidden_act[0] <= (hidden_sum[0] >= 5'sd0) ? 1'b1 : 1'b0;
                    hidden_act[1] <= (hidden_sum[1] >= 5'sd0) ? 1'b1 : 1'b0;
                    hidden_act[2] <= (hidden_sum[2] >= 5'sd0) ? 1'b1 : 1'b0;
                    hidden_act[3] <= (hidden_sum[3] >= 5'sd0) ? 1'b1 : 1'b0;
                    state <= COMPUTE_OUTPUT;
                end
                
                COMPUTE_OUTPUT: begin
                    classification <= decision;
                    state <= DONE;
                end
                
                DONE: begin
                    ready <= 1'b1;
                    state <= IDLE;  // Loop back for continuous monitoring
                end
                
                default: state <= IDLE;
            endcase
        end
    end
    
    // ========================================================================
    // OUTPUT PIN MAPPING
    // ========================================================================
    assign uo_out[0] = classification;           // 0=not ready, 1=ready to harvest
    assign uo_out[1] = ready;                    // Classification result ready
    assign uo_out[2] = (state == DONE);          // Processing complete indicator
    assign uo_out[3] = |inputs_binary;           // Any input active (sanity check)
    assign uo_out[7:4] = hidden_act;             // Debug: hidden layer state
    
endmodule
